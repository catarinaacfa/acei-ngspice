** Generated for: Eldo
** Generated on: Feb 27 10:58:28 2013
** Design library name: JoaoMelo
** Design cell name: Folded
** Design view name: Schematic

.OPTION TUNING=FAST
.OPTION AEX

.INC umc130.lib

.GLOBAL

.PARAM
+_vdd=3.3
+_wp5=2u
+_wp3=3u
+_wp1=2u
+_wp0=2u
+_wn7=2u
+_wn5=2u
+_wn3=2u 
+_wn2=2u
+_wn1=2u
+_nfp5=1
+_nfp3=1
+_nfp1=1
+_nfp0=1 
+_nfn7=1
+_nfn5=1
+_nfn3=1
+_nfn2=1
+_nfn1=1
+_lp1=360n
+_lp0=360n
+_ln7=360n
+_ln5=360n 
+_ln3=360n
+_ln1=360n


*********************************************************
** Library name: JoaoMelo
** Cell name: Folded
** View name: Schematic
.subckt Folded gnd ibias vdd vin vip vout
mnm7 net11 net11 gnd gnd N_HGLV_33_L130E w='_wn7/_nfn7' l=_ln7 as='_wn7/_nfn7<280e-9?(((78.4e-15+100e-9*(_wn7/_nfn7))+int((_nfn7-1)/2.0)*(78.4e-15+200e-9*(_wn7/_nfn7)))+(_nfn7/2-int(_nfn7/2)==0?78.4e-15+100e-9*(_wn7/_nfn7):0))/_nfn7:(((_wn7/_nfn7)*360e-9+int((_nfn7-1)/2.0)*((_wn7/_nfn7)*440e-9))+(_nfn7/2-int(_nfn7/2)==0?(_wn7/_nfn7)*360e-9:0))/_nfn7' ad='_wn7/_nfn7<280e-9?(int(_nfn7/2.0)*(78.4e-15+200e-9*(_wn7/_nfn7))+(_nfn7/2-int(_nfn7/2)!=0?78.4e-15+100e-9*(_wn7/_nfn7):0))/_nfn7:(int(_nfn7/2.0)*((_wn7/_nfn7)*440e-9)+(_nfn7/2-int(_nfn7/2)!=0?(_wn7/_nfn7)*360e-9:0))/_nfn7' ps='_wn7/_nfn7<280e-9?((1.32e-6+int((_nfn7-1)/2.0)*1.52e-6)+(_nfn7/2-int(_nfn7/2)==0?1.32e-6:0))/_nfn7:((2*(_wn7/_nfn7+360e-9)+int((_nfn7-1)/2.0)*(2*(_wn7/_nfn7+440e-9)))+(_nfn7/2-int(_nfn7/2)==0?2*(_wn7/_nfn7+360e-9):0))/_nfn7' pd='_wn7/_nfn7<280e-9?(int(_nfn7/2.0)*1.52e-6+(_nfn7/2-int(_nfn7/2)!=0?1.32e-6:0))/_nfn7:(int(_nfn7/2.0)*(2*(_wn7/_nfn7+440e-9))+(_nfn7/2-int(_nfn7/2)!=0?2*(_wn7/_nfn7+360e-9):0))/_nfn7' m='1*_nfn7'
mnm8 net15 net11 gnd gnd N_HGLV_33_L130E w='_wn7/_nfn7' l=_ln7 as='_wn7/_nfn7<280e-9?(((78.4e-15+100e-9*(_wn7/_nfn7))+int((_nfn7-1)/2.0)*(78.4e-15+200e-9*(_wn7/_nfn7)))+(_nfn7/2-int(_nfn7/2)==0?78.4e-15+100e-9*(_wn7/_nfn7):0))/_nfn7:(((_wn7/_nfn7)*360e-9+int((_nfn7-1)/2.0)*((_wn7/_nfn7)*440e-9))+(_nfn7/2-int(_nfn7/2)==0?(_wn7/_nfn7)*360e-9:0))/_nfn7' ad='_wn7/_nfn7<280e-9?(int(_nfn7/2.0)*(78.4e-15+200e-9*(_wn7/_nfn7))+(_nfn7/2-int(_nfn7/2)!=0?78.4e-15+100e-9*(_wn7/_nfn7):0))/_nfn7:(int(_nfn7/2.0)*((_wn7/_nfn7)*440e-9)+(_nfn7/2-int(_nfn7/2)!=0?(_wn7/_nfn7)*360e-9:0))/_nfn7' ps='_wn7/_nfn7<280e-9?((1.32e-6+int((_nfn7-1)/2.0)*1.52e-6)+(_nfn7/2-int(_nfn7/2)==0?1.32e-6:0))/_nfn7:((2*(_wn7/_nfn7+360e-9)+int((_nfn7-1)/2.0)*(2*(_wn7/_nfn7+440e-9)))+(_nfn7/2-int(_nfn7/2)==0?2*(_wn7/_nfn7+360e-9):0))/_nfn7' pd='_wn7/_nfn7<280e-9?(int(_nfn7/2.0)*1.52e-6+(_nfn7/2-int(_nfn7/2)!=0?1.32e-6:0))/_nfn7:(int(_nfn7/2.0)*(2*(_wn7/_nfn7+440e-9))+(_nfn7/2-int(_nfn7/2)!=0?2*(_wn7/_nfn7+360e-9):0))/_nfn7' m='1*_nfn7'
mnm2 net14 net27 gnd gnd N_HGLV_33_L130E w='_wn2/_nfn2' l=_ln1 as='_wn2/_nfn2<280e-9?(((78.4e-15+100e-9*(_wn2/_nfn2))+int((_nfn2-1)/2.0)*(78.4e-15+200e-9*(_wn2/_nfn2)))+(_nfn2/2-int(_nfn2/2)==0?78.4e-15+100e-9*(_wn2/_nfn2):0))/_nfn2:(((_wn2/_nfn2)*360e-9+int((_nfn2-1)/2.0)*((_wn2/_nfn2)*440e-9))+(_nfn2/2-int(_nfn2/2)==0?(_wn2/_nfn2)*360e-9:0))/_nfn2' ad='_wn2/_nfn2<280e-9?(int(_nfn2/2.0)*(78.4e-15+200e-9*(_wn2/_nfn2))+(_nfn2/2-int(_nfn2/2)!=0?78.4e-15+100e-9*(_wn2/_nfn2):0))/_nfn2:(int(_nfn2/2.0)*((_wn2/_nfn2)*440e-9)+(_nfn2/2-int(_nfn2/2)!=0?(_wn2/_nfn2)*360e-9:0))/_nfn2' ps='_wn2/_nfn2<280e-9?((1.32e-6+int((_nfn2-1)/2.0)*1.52e-6)+(_nfn2/2-int(_nfn2/2)==0?1.32e-6:0))/_nfn2:((2*(_wn2/_nfn2+360e-9)+int((_nfn2-1)/2.0)*(2*(_wn2/_nfn2+440e-9)))+(_nfn2/2-int(_nfn2/2)==0?2*(_wn2/_nfn2+360e-9):0))/_nfn2' pd='_wn2/_nfn2<280e-9?(int(_nfn2/2.0)*1.52e-6+(_nfn2/2-int(_nfn2/2)!=0?1.32e-6:0))/_nfn2:(int(_nfn2/2.0)*(2*(_wn2/_nfn2+440e-9))+(_nfn2/2-int(_nfn2/2)!=0?2*(_wn2/_nfn2+360e-9):0))/_nfn2' m='1*_nfn2'
mnm3 net0124 vip net14 net14 N_HGLV_33_L130E w='_wn3/_nfp3' l=_ln3 as='_wn3/_nfp3<280e-9?(((78.4e-15+100e-9*(_wn3/_nfp3))+int((_nfp3-1)/2.0)*(78.4e-15+200e-9*(_wn3/_nfp3)))+(_nfp3/2-int(_nfp3/2)==0?78.4e-15+100e-9*(_wn3/_nfp3):0))/_nfp3:(((_wn3/_nfp3)*360e-9+int((_nfp3-1)/2.0)*((_wn3/_nfp3)*440e-9))+(_nfp3/2-int(_nfp3/2)==0?(_wn3/_nfp3)*360e-9:0))/_nfp3' ad='_wn3/_nfp3<280e-9?(int(_nfp3/2.0)*(78.4e-15+200e-9*(_wn3/_nfp3))+(_nfp3/2-int(_nfp3/2)!=0?78.4e-15+100e-9*(_wn3/_nfp3):0))/_nfp3:(int(_nfp3/2.0)*((_wn3/_nfp3)*440e-9)+(_nfp3/2-int(_nfp3/2)!=0?(_wn3/_nfp3)*360e-9:0))/_nfp3' ps='_wn3/_nfp3<280e-9?((1.32e-6+int((_nfp3-1)/2.0)*1.52e-6)+(_nfp3/2-int(_nfp3/2)==0?1.32e-6:0))/_nfp3:((2*(_wn3/_nfp3+360e-9)+int((_nfp3-1)/2.0)*(2*(_wn3/_nfp3+440e-9)))+(_nfp3/2-int(_nfp3/2)==0?2*(_wn3/_nfp3+360e-9):0))/_nfp3' pd='_wn3/_nfp3<280e-9?(int(_nfp3/2.0)*1.52e-6+(_nfp3/2-int(_nfp3/2)!=0?1.32e-6:0))/_nfp3:(int(_nfp3/2.0)*(2*(_wn3/_nfp3+440e-9))+(_nfp3/2-int(_nfp3/2)!=0?2*(_wn3/_nfp3+360e-9):0))/_nfp3' m='1*_nfp3'
mnm4 net0128 vin net14 net14 N_HGLV_33_L130E w='_wn3/_nfn3' l=_ln3 as='_wn3/_nfn3<280e-9?(((78.4e-15+100e-9*(_wn3/_nfn3))+int((_nfn3-1)/2.0)*(78.4e-15+200e-9*(_wn3/_nfn3)))+(_nfn3/2-int(_nfn3/2)==0?78.4e-15+100e-9*(_wn3/_nfn3):0))/_nfn3:(((_wn3/_nfn3)*360e-9+int((_nfn3-1)/2.0)*((_wn3/_nfn3)*440e-9))+(_nfn3/2-int(_nfn3/2)==0?(_wn3/_nfn3)*360e-9:0))/_nfn3' ad='_wn3/_nfn3<280e-9?(int(_nfn3/2.0)*(78.4e-15+200e-9*(_wn3/_nfn3))+(_nfn3/2-int(_nfn3/2)!=0?78.4e-15+100e-9*(_wn3/_nfn3):0))/_nfn3:(int(_nfn3/2.0)*((_wn3/_nfn3)*440e-9)+(_nfn3/2-int(_nfn3/2)!=0?(_wn3/_nfn3)*360e-9:0))/_nfn3' ps='_wn3/_nfn3<280e-9?((1.32e-6+int((_nfn3-1)/2.0)*1.52e-6)+(_nfn3/2-int(_nfn3/2)==0?1.32e-6:0))/_nfn3:((2*(_wn3/_nfn3+360e-9)+int((_nfn3-1)/2.0)*(2*(_wn3/_nfn3+440e-9)))+(_nfn3/2-int(_nfn3/2)==0?2*(_wn3/_nfn3+360e-9):0))/_nfn3' pd='_wn3/_nfn3<280e-9?(int(_nfn3/2.0)*1.52e-6+(_nfn3/2-int(_nfn3/2)!=0?1.32e-6:0))/_nfn3:(int(_nfn3/2.0)*(2*(_wn3/_nfn3+440e-9))+(_nfn3/2-int(_nfn3/2)!=0?2*(_wn3/_nfn3+360e-9):0))/_nfn3' m='1*_nfn3'
mnm6 vout net31 net15 net15 N_HGLV_33_L130E w='_wn5/_nfn5' l=_ln5 as='_wn5/_nfn5<280e-9?(((78.4e-15+100e-9*(_wn5/_nfn5))+int((_nfn5-1)/2.0)*(78.4e-15+200e-9*(_wn5/_nfn5)))+(_nfn5/2-int(_nfn5/2)==0?78.4e-15+100e-9*(_wn5/_nfn5):0))/_nfn5:(((_wn5/_nfn5)*360e-9+int((_nfn5-1)/2.0)*((_wn5/_nfn5)*440e-9))+(_nfn5/2-int(_nfn5/2)==0?(_wn5/_nfn5)*360e-9:0))/_nfn5' ad='_wn5/_nfn5<280e-9?(int(_nfn5/2.0)*(78.4e-15+200e-9*(_wn5/_nfn5))+(_nfn5/2-int(_nfn5/2)!=0?78.4e-15+100e-9*(_wn5/_nfn5):0))/_nfn5:(int(_nfn5/2.0)*((_wn5/_nfn5)*440e-9)+(_nfn5/2-int(_nfn5/2)!=0?(_wn5/_nfn5)*360e-9:0))/_nfn5' ps='_wn5/_nfn5<280e-9?((1.32e-6+int((_nfn5-1)/2.0)*1.52e-6)+(_nfn5/2-int(_nfn5/2)==0?1.32e-6:0))/_nfn5:((2*(_wn5/_nfn5+360e-9)+int((_nfn5-1)/2.0)*(2*(_wn5/_nfn5+440e-9)))+(_nfn5/2-int(_nfn5/2)==0?2*(_wn5/_nfn5+360e-9):0))/_nfn5' pd='_wn5/_nfn5<280e-9?(int(_nfn5/2.0)*1.52e-6+(_nfn5/2-int(_nfn5/2)!=0?1.32e-6:0))/_nfn5:(int(_nfn5/2.0)*(2*(_wn5/_nfn5+440e-9))+(_nfn5/2-int(_nfn5/2)!=0?2*(_wn5/_nfn5+360e-9):0))/_nfn5' m='1*_nfn5'
mnm5 net31 net31 net11 net11 N_HGLV_33_L130E w='_wn5/_nfn5' l=_ln5 as='_wn5/_nfn5<280e-9?(((78.4e-15+100e-9*(_wn5/_nfn5))+int((_nfn5-1)/2.0)*(78.4e-15+200e-9*(_wn5/_nfn5)))+(_nfn5/2-int(_nfn5/2)==0?78.4e-15+100e-9*(_wn5/_nfn5):0))/_nfn5:(((_wn5/_nfn5)*360e-9+int((_nfn5-1)/2.0)*((_wn5/_nfn5)*440e-9))+(_nfn5/2-int(_nfn5/2)==0?(_wn5/_nfn5)*360e-9:0))/_nfn5' ad='_wn5/_nfn5<280e-9?(int(_nfn5/2.0)*(78.4e-15+200e-9*(_wn5/_nfn5))+(_nfn5/2-int(_nfn5/2)!=0?78.4e-15+100e-9*(_wn5/_nfn5):0))/_nfn5:(int(_nfn5/2.0)*((_wn5/_nfn5)*440e-9)+(_nfn5/2-int(_nfn5/2)!=0?(_wn5/_nfn5)*360e-9:0))/_nfn5' ps='_wn5/_nfn5<280e-9?((1.32e-6+int((_nfn5-1)/2.0)*1.52e-6)+(_nfn5/2-int(_nfn5/2)==0?1.32e-6:0))/_nfn5:((2*(_wn5/_nfn5+360e-9)+int((_nfn5-1)/2.0)*(2*(_wn5/_nfn5+440e-9)))+(_nfn5/2-int(_nfn5/2)==0?2*(_wn5/_nfn5+360e-9):0))/_nfn5' pd='_wn5/_nfn5<280e-9?(int(_nfn5/2.0)*1.52e-6+(_nfn5/2-int(_nfn5/2)!=0?1.32e-6:0))/_nfn5:(int(_nfn5/2.0)*(2*(_wn5/_nfn5+440e-9))+(_nfn5/2-int(_nfn5/2)!=0?2*(_wn5/_nfn5+360e-9):0))/_nfn5' m='1*_nfn5'
mnm1 net27 net27 gnd gnd N_HGLV_33_L130E w='_wn1/_nfn1' l=_ln1 as='_wn1/_nfn1<280e-9?(((78.4e-15+100e-9*(_wn1/_nfn1))+int((_nfn1-1)/2.0)*(78.4e-15+200e-9*(_wn1/_nfn1)))+(_nfn1/2-int(_nfn1/2)==0?78.4e-15+100e-9*(_wn1/_nfn1):0))/_nfn1:(((_wn1/_nfn1)*360e-9+int((_nfn1-1)/2.0)*((_wn1/_nfn1)*440e-9))+(_nfn1/2-int(_nfn1/2)==0?(_wn1/_nfn1)*360e-9:0))/_nfn1' ad='_wn1/_nfn1<280e-9?(int(_nfn1/2.0)*(78.4e-15+200e-9*(_wn1/_nfn1))+(_nfn1/2-int(_nfn1/2)!=0?78.4e-15+100e-9*(_wn1/_nfn1):0))/_nfn1:(int(_nfn1/2.0)*((_wn1/_nfn1)*440e-9)+(_nfn1/2-int(_nfn1/2)!=0?(_wn1/_nfn1)*360e-9:0))/_nfn1' ps='_wn1/_nfn1<280e-9?((1.32e-6+int((_nfn1-1)/2.0)*1.52e-6)+(_nfn1/2-int(_nfn1/2)==0?1.32e-6:0))/_nfn1:((2*(_wn1/_nfn1+360e-9)+int((_nfn1-1)/2.0)*(2*(_wn1/_nfn1+440e-9)))+(_nfn1/2-int(_nfn1/2)==0?2*(_wn1/_nfn1+360e-9):0))/_nfn1' pd='_wn1/_nfn1<280e-9?(int(_nfn1/2.0)*1.52e-6+(_nfn1/2-int(_nfn1/2)!=0?1.32e-6:0))/_nfn1:(int(_nfn1/2.0)*(2*(_wn1/_nfn1+440e-9))+(_nfn1/2-int(_nfn1/2)!=0?2*(_wn1/_nfn1+360e-9):0))/_nfn1' m='1*_nfn1'
mpm4 net0128 net56 vdd vdd P_HGLV_33_L130E w='_wp3/_nfp3' l=_lp0 as='_wp3/_nfp3<280e-9?(((78.4e-15+100e-9*(_wp3/_nfp3))+int((_nfp3-1)/2.0)*(78.4e-15+200e-9*(_wp3/_nfp3)))+(_nfp3/2-int(_nfp3/2)==0?78.4e-15+100e-9*(_wp3/_nfp3):0))/_nfp3:(((_wp3/_nfp3)*360e-9+int((_nfp3-1)/2.0)*((_wp3/_nfp3)*440e-9))+(_nfp3/2-int(_nfp3/2)==0?(_wp3/_nfp3)*360e-9:0))/_nfp3' ad='_wp3/_nfp3<280e-9?(int(_nfp3/2.0)*(78.4e-15+200e-9*(_wp3/_nfp3))+(_nfp3/2-int(_nfp3/2)!=0?78.4e-15+100e-9*(_wp3/_nfp3):0))/_nfp3:(int(_nfp3/2.0)*((_wp3/_nfp3)*440e-9)+(_nfp3/2-int(_nfp3/2)!=0?(_wp3/_nfp3)*360e-9:0))/_nfp3' ps='_wp3/_nfp3<280e-9?((1.32e-6+int((_nfp3-1)/2.0)*1.52e-6)+(_nfp3/2-int(_nfp3/2)==0?1.32e-6:0))/_nfp3:((2*(_wp3/_nfp3+360e-9)+int((_nfp3-1)/2.0)*(2*(_wp3/_nfp3+440e-9)))+(_nfp3/2-int(_nfp3/2)==0?2*(_wp3/_nfp3+360e-9):0))/_nfp3' pd='_wp3/_nfp3<280e-9?(int(_nfp3/2.0)*1.52e-6+(_nfp3/2-int(_nfp3/2)!=0?1.32e-6:0))/_nfp3:(int(_nfp3/2.0)*(2*(_wp3/_nfp3+440e-9))+(_nfp3/2-int(_nfp3/2)!=0?2*(_wp3/_nfp3+360e-9):0))/_nfp3' m='1*_nfp3'
mpm3 net0124 net56 vdd vdd P_HGLV_33_L130E w='_wp3/_nfp3' l=_lp0 as='_wp3/_nfp3<280e-9?(((78.4e-15+100e-9*(_wp3/_nfp3))+int((_nfp3-1)/2.0)*(78.4e-15+200e-9*(_wp3/_nfp3)))+(_nfp3/2-int(_nfp3/2)==0?78.4e-15+100e-9*(_wp3/_nfp3):0))/_nfp3:(((_wp3/_nfp3)*360e-9+int((_nfp3-1)/2.0)*((_wp3/_nfp3)*440e-9))+(_nfp3/2-int(_nfp3/2)==0?(_wp3/_nfp3)*360e-9:0))/_nfp3' ad='_wp3/_nfp3<280e-9?(int(_nfp3/2.0)*(78.4e-15+200e-9*(_wp3/_nfp3))+(_nfp3/2-int(_nfp3/2)!=0?78.4e-15+100e-9*(_wp3/_nfp3):0))/_nfp3:(int(_nfp3/2.0)*((_wp3/_nfp3)*440e-9)+(_nfp3/2-int(_nfp3/2)!=0?(_wp3/_nfp3)*360e-9:0))/_nfp3' ps='_wp3/_nfp3<280e-9?((1.32e-6+int((_nfp3-1)/2.0)*1.52e-6)+(_nfp3/2-int(_nfp3/2)==0?1.32e-6:0))/_nfp3:((2*(_wp3/_nfp3+360e-9)+int((_nfp3-1)/2.0)*(2*(_wp3/_nfp3+440e-9)))+(_nfp3/2-int(_nfp3/2)==0?2*(_wp3/_nfp3+360e-9):0))/_nfp3' pd='_wp3/_nfp3<280e-9?(int(_nfp3/2.0)*1.52e-6+(_nfp3/2-int(_nfp3/2)!=0?1.32e-6:0))/_nfp3:(int(_nfp3/2.0)*(2*(_wp3/_nfp3+440e-9))+(_nfp3/2-int(_nfp3/2)!=0?2*(_wp3/_nfp3+360e-9):0))/_nfp3' m='1*_nfp3'
mpm6 vout net27 net0128 net0128 P_HGLV_33_L130E w='_wp5/_nfp5' l=_lp1 as='_wp5/_nfp5<280e-9?(((78.4e-15+100e-9*(_wp5/_nfp5))+int((_nfp5-1)/2.0)*(78.4e-15+200e-9*(_wp5/_nfp5)))+(_nfp5/2-int(_nfp5/2)==0?78.4e-15+100e-9*(_wp5/_nfp5):0))/_nfp5:(((_wp5/_nfp5)*360e-9+int((_nfp5-1)/2.0)*((_wp5/_nfp5)*440e-9))+(_nfp5/2-int(_nfp5/2)==0?(_wp5/_nfp5)*360e-9:0))/_nfp5' ad='_wp5/_nfp5<280e-9?(int(_nfp5/2.0)*(78.4e-15+200e-9*(_wp5/_nfp5))+(_nfp5/2-int(_nfp5/2)!=0?78.4e-15+100e-9*(_wp5/_nfp5):0))/_nfp5:(int(_nfp5/2.0)*((_wp5/_nfp5)*440e-9)+(_nfp5/2-int(_nfp5/2)!=0?(_wp5/_nfp5)*360e-9:0))/_nfp5' ps='_wp5/_nfp5<280e-9?((1.32e-6+int((_nfp5-1)/2.0)*1.52e-6)+(_nfp5/2-int(_nfp5/2)==0?1.32e-6:0))/_nfp5:((2*(_wp5/_nfp5+360e-9)+int((_nfp5-1)/2.0)*(2*(_wp5/_nfp5+440e-9)))+(_nfp5/2-int(_nfp5/2)==0?2*(_wp5/_nfp5+360e-9):0))/_nfp5' pd='_wp5/_nfp5<280e-9?(int(_nfp5/2.0)*1.52e-6+(_nfp5/2-int(_nfp5/2)!=0?1.32e-6:0))/_nfp5:(int(_nfp5/2.0)*(2*(_wp5/_nfp5+440e-9))+(_nfp5/2-int(_nfp5/2)!=0?2*(_wp5/_nfp5+360e-9):0))/_nfp5' m='1*_nfp5'
mpm0 net56 net56 ibias ibias P_HGLV_33_L130E w='_wp0/_nfp0' l=_lp0 as='_wp0/_nfp0<280e-9?(((78.4e-15+100e-9*(_wp0/_nfp0))+int((_nfp0-1)/2.0)*(78.4e-15+200e-9*(_wp0/_nfp0)))+(_nfp0/2-int(_nfp0/2)==0?78.4e-15+100e-9*(_wp0/_nfp0):0))/_nfp0:(((_wp0/_nfp0)*360e-9+int((_nfp0-1)/2.0)*((_wp0/_nfp0)*440e-9))+(_nfp0/2-int(_nfp0/2)==0?(_wp0/_nfp0)*360e-9:0))/_nfp0' ad='_wp0/_nfp0<280e-9?(int(_nfp0/2.0)*(78.4e-15+200e-9*(_wp0/_nfp0))+(_nfp0/2-int(_nfp0/2)!=0?78.4e-15+100e-9*(_wp0/_nfp0):0))/_nfp0:(int(_nfp0/2.0)*((_wp0/_nfp0)*440e-9)+(_nfp0/2-int(_nfp0/2)!=0?(_wp0/_nfp0)*360e-9:0))/_nfp0' ps='_wp0/_nfp0<280e-9?((1.32e-6+int((_nfp0-1)/2.0)*1.52e-6)+(_nfp0/2-int(_nfp0/2)==0?1.32e-6:0))/_nfp0:((2*(_wp0/_nfp0+360e-9)+int((_nfp0-1)/2.0)*(2*(_wp0/_nfp0+440e-9)))+(_nfp0/2-int(_nfp0/2)==0?2*(_wp0/_nfp0+360e-9):0))/_nfp0' pd='_wp0/_nfp0<280e-9?(int(_nfp0/2.0)*1.52e-6+(_nfp0/2-int(_nfp0/2)!=0?1.32e-6:0))/_nfp0:(int(_nfp0/2.0)*(2*(_wp0/_nfp0+440e-9))+(_nfp0/2-int(_nfp0/2)!=0?2*(_wp0/_nfp0+360e-9):0))/_nfp0' m='1*_nfp0'
mpm5 net31 net27 net0124 net0124 P_HGLV_33_L130E w='_wp5/_nfp5' l=_lp1 as='_wp5/_nfp5<280e-9?(((78.4e-15+100e-9*(_wp5/_nfp5))+int((_nfp5-1)/2.0)*(78.4e-15+200e-9*(_wp5/_nfp5)))+(_nfp5/2-int(_nfp5/2)==0?78.4e-15+100e-9*(_wp5/_nfp5):0))/_nfp5:(((_wp5/_nfp5)*360e-9+int((_nfp5-1)/2.0)*((_wp5/_nfp5)*440e-9))+(_nfp5/2-int(_nfp5/2)==0?(_wp5/_nfp5)*360e-9:0))/_nfp5' ad='_wp5/_nfp5<280e-9?(int(_nfp5/2.0)*(78.4e-15+200e-9*(_wp5/_nfp5))+(_nfp5/2-int(_nfp5/2)!=0?78.4e-15+100e-9*(_wp5/_nfp5):0))/_nfp5:(int(_nfp5/2.0)*((_wp5/_nfp5)*440e-9)+(_nfp5/2-int(_nfp5/2)!=0?(_wp5/_nfp5)*360e-9:0))/_nfp5' ps='_wp5/_nfp5<280e-9?((1.32e-6+int((_nfp5-1)/2.0)*1.52e-6)+(_nfp5/2-int(_nfp5/2)==0?1.32e-6:0))/_nfp5:((2*(_wp5/_nfp5+360e-9)+int((_nfp5-1)/2.0)*(2*(_wp5/_nfp5+440e-9)))+(_nfp5/2-int(_nfp5/2)==0?2*(_wp5/_nfp5+360e-9):0))/_nfp5' pd='_wp5/_nfp5<280e-9?(int(_nfp5/2.0)*1.52e-6+(_nfp5/2-int(_nfp5/2)!=0?1.32e-6:0))/_nfp5:(int(_nfp5/2.0)*(2*(_wp5/_nfp5+440e-9))+(_nfp5/2-int(_nfp5/2)!=0?2*(_wp5/_nfp5+360e-9):0))/_nfp5' m='1*_nfp5'
mpm1 net27 net27 net56 net56 P_HGLV_33_L130E w='_wp1/_nfp1' l=_lp1 as='_wp1/_nfp1<280e-9?(((78.4e-15+100e-9*(_wp1/_nfp1))+int((_nfp1-1)/2.0)*(78.4e-15+200e-9*(_wp1/_nfp1)))+(_nfp1/2-int(_nfp1/2)==0?78.4e-15+100e-9*(_wp1/_nfp1):0))/_nfp1:(((_wp1/_nfp1)*360e-9+int((_nfp1-1)/2.0)*((_wp1/_nfp1)*440e-9))+(_nfp1/2-int(_nfp1/2)==0?(_wp1/_nfp1)*360e-9:0))/_nfp1' ad='_wp1/_nfp1<280e-9?(int(_nfp1/2.0)*(78.4e-15+200e-9*(_wp1/_nfp1))+(_nfp1/2-int(_nfp1/2)!=0?78.4e-15+100e-9*(_wp1/_nfp1):0))/_nfp1:(int(_nfp1/2.0)*((_wp1/_nfp1)*440e-9)+(_nfp1/2-int(_nfp1/2)!=0?(_wp1/_nfp1)*360e-9:0))/_nfp1' ps='_wp1/_nfp1<280e-9?((1.32e-6+int((_nfp1-1)/2.0)*1.52e-6)+(_nfp1/2-int(_nfp1/2)==0?1.32e-6:0))/_nfp1:((2*(_wp1/_nfp1+360e-9)+int((_nfp1-1)/2.0)*(2*(_wp1/_nfp1+440e-9)))+(_nfp1/2-int(_nfp1/2)==0?2*(_wp1/_nfp1+360e-9):0))/_nfp1' pd='_wp1/_nfp1<280e-9?(int(_nfp1/2.0)*1.52e-6+(_nfp1/2-int(_nfp1/2)!=0?1.32e-6:0))/_nfp1:(int(_nfp1/2.0)*(2*(_wp1/_nfp1+440e-9))+(_nfp1/2-int(_nfp1/2)!=0?2*(_wp1/_nfp1+360e-9):0))/_nfp1' m='1*_nfp1'
.ends
*********************************************************

*********************************************************
** Library name: JoaoMelo
** Cell name: Testbench
** View name: Schematic
xi10 0 net15 vddnet vin vip vout Folded
c0 vout 0 10e-12
v2 vin 0 DC=1.65	
v1 vip 0 DC=1.65 AC 1
v0 vddnet 0 DC=_vdd
i1 vddnet net15 DC=100u

xi11 0 net16 vddd vinn vipp voutt Folded
c1 voutt 0 10e-12
v5 vipp 0 DC=1.65
v4 vinn 0 DC=1.65
v3 vddd 0 DC=_vdd AC 1
i2 vddd net16 DC=100u
*********************************************************

*********** Analysis ***************************
.TEMP 25.0
*.AC DEC 200 1 1G 
.OPTION BRIEF=0
************************************************


.control

set units = degrees

AC DEC 200 1 1G

meas AC GDC FIND vdb(vout) at=1
meas AC GBW WHEN vdb(vout)=0
meas AC PM FIND vp(vout) WHEN vdb(vout)=0
meas AC GPS FIND vdb(voutt) at=1

let PSRR = GDC-GPS
print PSRR

let ids = @m.xi10.mpm6[id]
print ids

let SR = (ids/10E-12)*1E-6
print SR

quit


.endc


.END
